//----------------------------------------------------------------------
// seizure_detection_tb.sv
// Testbench for epileptic seizure detection system
//----------------------------------------------------------------------

module seizure_detection_tb;
    // Parameters
    localparam DATA_WIDTH = 16;
    localparam FEATURE_COUNT = 178;
    localparam CLK_PERIOD = 10; // 10ns (100MHz)
    localparam TEST_VECTORS = 10;
    
    // Signals
    logic clk;
    logic rst_n;
    logic data_valid;
    logic [DATA_WIDTH-1:0] eeg_data [FEATURE_COUNT-1:0];
    logic system_ready;
    logic result_valid;
    logic seizure_detected;
    logic [DATA_WIDTH-1:0] detection_confidence;
    logic [1:0] system_status;
    
    // Test vector storage
    logic [DATA_WIDTH-1:0] test_vectors [TEST_VECTORS-1:0][FEATURE_COUNT-1:0];
    logic expected_results [TEST_VECTORS-1:0];
    
    // Statistics
    integer correct_classifications;
    integer total_tests;
    real accuracy;
    
    // DUT instantiation
    seizure_detection_system #(
        .DATA_WIDTH(DATA_WIDTH),
        .FEATURE_COUNT(FEATURE_COUNT)
    ) dut (
        .clk(clk),
        .rst_n(rst_n),
        .data_valid(data_valid),
        .eeg_data(eeg_data),
        .system_ready(system_ready),
        .result_valid(result_valid),
        .seizure_detected(seizure_detected),
        .detection_confidence(detection_confidence),
        .system_status(system_status)
    );
    
    // Clock generation
    initial begin
        clk = 0;
        forever #(CLK_PERIOD/2) clk = ~clk;
    end
    
    // Reset generation
    initial begin
        rst_n = 0;
        #(CLK_PERIOD*5) rst_n = 1;
    end
    
    // Load test vectors
    initial begin
        // In practice, you would load these from a file generated by your Python script
        // For now, we'll create synthetic test data
        for (int i = 0; i < TEST_VECTORS; i++) begin
            // Even test vectors are seizure cases (class 1)
            // Odd test vectors are non-seizure cases (classes 2-5)
            expected_results[i] = (i % 2 == 0);
            
            for (int j = 0; j < FEATURE_COUNT; j++) begin
                if (expected_results[i]) 
                    // Seizure pattern
                    test_vectors[i][j] = 16'h0100 + ((i*j) & 16'h00FF);
                else
                    // Non-seizure pattern
                    test_vectors[i][j] = 16'h0200 + ((i*j) & 16'h00FF);
            end
        end
        
        correct_classifications = 0;
        total_tests = 0;
    end
    
    // Test process
    initial begin
        data_valid = 0;
        
        // Wait for reset and initialization
        wait(rst_n);
        repeat(5) @(posedge clk);
        
        // Run through test vectors
        for (int i = 0; i < TEST_VECTORS; i++) begin
            $display("Running test vector %0d...", i);
            
            // Wait until system is ready
            wait(system_ready);
            @(posedge clk);
            
            // Load test vector
            for (int j = 0; j < FEATURE_COUNT; j++) begin
                eeg_data[j] = test_vectors[i][j];
            end
            
            // Signal data is valid
            data_valid = 1;
            @(posedge clk);
            data_valid = 0;
            
            // Wait for result
            wait(result_valid);
            @(posedge clk);
            
            // Check result
            total_tests++;
            if (seizure_detected == expected_results[i]) begin
                correct_classifications++;
                $display("Test %0d: PASSED - Expected: %s, Got: %s, Confidence: %f", 
                       i, 
                       expected_results[i] ? "Seizure" : "Non-seizure",
                       seizure_detected ? "Seizure" : "Non-seizure",
                       real'(detection_confidence) / 256.0);
            end else begin
                $display("Test %0d: FAILED - Expected: %s, Got: %s, Confidence: %f", 
                       i, 
                       expected_results[i] ? "Seizure" : "Non-seizure",
                       seizure_detected ? "Seizure" : "Non-seizure",
                       real'(detection_confidence) / 256.0);
            end
            
            // Wait between tests
            repeat(10) @(posedge clk);
        end
        
        // Calculate and display accuracy
        accuracy = 100.0 * real'(correct_classifications) / real'(total_tests);
        
        $display("\n===== Test Results =====");
        $display("Total tests: %0d", total_tests);
        $display("Correct classifications: %0d", correct_classifications);
        $display("Accuracy: %.2f%%", accuracy);
        $display("=======================\n");
        
        // End simulation
        #100 $finish;
    end
    
    // Monitor key signals
    initial begin
        $monitor("Time: %t, State: %s, Ready: %b, Valid: %b", 
                $time, 
                system_status == 0 ? "IDLE" : 
                system_status == 1 ? "PROCESSING" : 
                system_status == 2 ? "RESULT_READY" : "ERROR",
                system_ready, 
                result_valid);
    end

endmodule